`ifndef CFS_MD_PKG_SV
    `define CFS_MD_PKG_SV

    // `include "uvm_macros.svh"
    `include "cfs_md_if.sv"

    package cfs_md_pkg;
        // import uvm_pkg::*;

    endpackage
`endif
